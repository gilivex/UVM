// header - package file to include the env and test
package my_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "my_transaction.sv"
	`include "my_sequencer.sv"
	`include "my_sequence.sv"	
	`include "my_driver.sv"
	`include "my_agent.sv"
	`include "my_env.sv"
	`include "random_test.sv"
	
endpackage